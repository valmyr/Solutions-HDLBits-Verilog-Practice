module step_One( output one );
    assign one = 1;
endmodule