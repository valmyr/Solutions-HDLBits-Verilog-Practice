/*
We're going to start with a small bit of HDL to get familiar with the interface used by HDLBits. Here's the description of the circuit you need to build for this exercise:

Build a circuit with no inputs and one output. That output should always drive 1 (or logic high).


Expected solution length: Around 1 line.

*/

module testBenchStep_One();
  logic one;
  step_One oneInsta(one);
  initial begin
    $monitor("%b",one);
  end
endmodule